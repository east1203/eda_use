module add (input a,b,c,d ,output sum1,sum2);

assign sum1 = a+b+c+d;
assign sum2 =(a+b) + (c+d);

endmodule
